module Baud_Rate_Generator ();


  
endmodule
